module main

pub struct Config {
pub:
    title string = 'My Docs'
}
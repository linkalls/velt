module main

pub struct Config {
pub:
    title string = 'My Blog'
    theme string = 'blog'
}